// clkmux_cv.v

// Generated using ACDS version 14.1 186 at 2014.12.20.10:36:39

`timescale 1 ps / 1 ps
module clkmux_cv (
		input  wire       inclk2x,   //  altclkctrl_input.inclk2x
		input  wire       inclk1x,   //                  .inclk1x
		input  wire       inclk0x,   //                  .inclk0x
		input  wire [1:0] clkselect, //                  .clkselect
		output wire       outclk     // altclkctrl_output.outclk
	);

	clkmux_cv_altclkctrl_0 altclkctrl_0 (
		.inclk2x   (inclk2x),   //  altclkctrl_input.inclk2x
		.inclk1x   (inclk1x),   //                  .inclk1x
		.inclk0x   (inclk0x),   //                  .inclk0x
		.clkselect (clkselect), //                  .clkselect
		.outclk    (outclk)     // altclkctrl_output.outclk
	);

endmodule
