// megafunction wizard: %ALTASMI_PARALLEL%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTASMI_PARALLEL 

// ============================================================
// File Name: ASMI.v
// Megafunction Name(s):
// 			ALTASMI_PARALLEL
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 14.0.1 Build 205 08/13/2014 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, the Altera Quartus II License Agreement,
//the Altera MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Altera and sold by Altera or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.

module ASMI (
	addr,
	bulk_erase,
	clkin,
	datain,
	rden,
	read,
	read_sid,
	reset,
	sector_erase,
	sector_protect,
	shift_bytes,
	wren,
	write,
	busy,
	data_valid,
	dataout,
	epcs_id,
	illegal_erase,
	illegal_write)/* synthesis synthesis_clearbox = 1 */;

	input	[23:0]  addr;
	input	  bulk_erase;
	input	  clkin;
	input	[7:0]  datain;
	input	  rden;
	input	  read;
	input	  read_sid;
	input	  reset;
	input	  sector_erase;
	input	  sector_protect;
	input	  shift_bytes;
	input	  wren;
	input	  write;
	output	  busy;
	output	  data_valid;
	output	[7:0]  dataout;
	output	[7:0]  epcs_id;
	output	  illegal_erase;
	output	  illegal_write;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: DATA_WIDTH STRING "STANDARD"
// Retrieval info: CONSTANT: ENABLE_SIM STRING "FALSE"
// Retrieval info: CONSTANT: EPCS_TYPE STRING "EPCS16"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altasmi_parallel"
// Retrieval info: CONSTANT: PAGE_SIZE NUMERIC "256"
// Retrieval info: CONSTANT: PORT_BULK_ERASE STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_DIE_ERASE STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_EN4B_ADDR STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_EX4B_ADDR STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_FAST_READ STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_ILLEGAL_ERASE STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_ILLEGAL_WRITE STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_RDID_OUT STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_READ_ADDRESS STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_READ_DUMMYCLK STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_READ_RDID STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_READ_SID STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_READ_STATUS STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SECTOR_ERASE STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_SECTOR_PROTECT STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_SHIFT_BYTES STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_WREN STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_WRITE STRING "PORT_USED"
// Retrieval info: CONSTANT: USE_ASMIBLOCK STRING "ON"
// Retrieval info: CONSTANT: USE_EAB STRING "ON"
// Retrieval info: CONSTANT: WRITE_DUMMY_CLK NUMERIC "0"
// Retrieval info: USED_PORT: addr 0 0 24 0 INPUT NODEFVAL "addr[23..0]"
// Retrieval info: CONNECT: @addr 0 0 24 0 addr 0 0 24 0
// Retrieval info: USED_PORT: bulk_erase 0 0 0 0 INPUT NODEFVAL "bulk_erase"
// Retrieval info: CONNECT: @bulk_erase 0 0 0 0 bulk_erase 0 0 0 0
// Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
// Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
// Retrieval info: USED_PORT: clkin 0 0 0 0 INPUT NODEFVAL "clkin"
// Retrieval info: CONNECT: @clkin 0 0 0 0 clkin 0 0 0 0
// Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
// Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
// Retrieval info: USED_PORT: datain 0 0 8 0 INPUT NODEFVAL "datain[7..0]"
// Retrieval info: CONNECT: @datain 0 0 8 0 datain 0 0 8 0
// Retrieval info: USED_PORT: dataout 0 0 8 0 OUTPUT NODEFVAL "dataout[7..0]"
// Retrieval info: CONNECT: dataout 0 0 8 0 @dataout 0 0 8 0
// Retrieval info: USED_PORT: epcs_id 0 0 8 0 OUTPUT NODEFVAL "epcs_id[7..0]"
// Retrieval info: CONNECT: epcs_id 0 0 8 0 @epcs_id 0 0 8 0
// Retrieval info: USED_PORT: illegal_erase 0 0 0 0 OUTPUT NODEFVAL "illegal_erase"
// Retrieval info: CONNECT: illegal_erase 0 0 0 0 @illegal_erase 0 0 0 0
// Retrieval info: USED_PORT: illegal_write 0 0 0 0 OUTPUT NODEFVAL "illegal_write"
// Retrieval info: CONNECT: illegal_write 0 0 0 0 @illegal_write 0 0 0 0
// Retrieval info: USED_PORT: rden 0 0 0 0 INPUT NODEFVAL "rden"
// Retrieval info: CONNECT: @rden 0 0 0 0 rden 0 0 0 0
// Retrieval info: USED_PORT: read 0 0 0 0 INPUT NODEFVAL "read"
// Retrieval info: CONNECT: @read 0 0 0 0 read 0 0 0 0
// Retrieval info: USED_PORT: read_sid 0 0 0 0 INPUT NODEFVAL "read_sid"
// Retrieval info: CONNECT: @read_sid 0 0 0 0 read_sid 0 0 0 0
// Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
// Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
// Retrieval info: USED_PORT: sector_erase 0 0 0 0 INPUT NODEFVAL "sector_erase"
// Retrieval info: CONNECT: @sector_erase 0 0 0 0 sector_erase 0 0 0 0
// Retrieval info: USED_PORT: sector_protect 0 0 0 0 INPUT NODEFVAL "sector_protect"
// Retrieval info: CONNECT: @sector_protect 0 0 0 0 sector_protect 0 0 0 0
// Retrieval info: USED_PORT: shift_bytes 0 0 0 0 INPUT NODEFVAL "shift_bytes"
// Retrieval info: CONNECT: @shift_bytes 0 0 0 0 shift_bytes 0 0 0 0
// Retrieval info: USED_PORT: wren 0 0 0 0 INPUT NODEFVAL "wren"
// Retrieval info: CONNECT: @wren 0 0 0 0 wren 0 0 0 0
// Retrieval info: USED_PORT: write 0 0 0 0 INPUT NODEFVAL "write"
// Retrieval info: CONNECT: @write 0 0 0 0 write 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL ASMI.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ASMI.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ASMI.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ASMI_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ASMI_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ASMI.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ASMI.cmp TRUE TRUE
